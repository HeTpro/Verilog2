module nombre(a, b, c);
  input s

endmodule
